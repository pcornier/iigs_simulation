// 
// Apple ][ track read/write interface to MiST
//
// Based on the work of
// Copyright (c) 2016 Sorgelig
//
// This source file is free software: you can redistribute it and/or modify
// it under the terms of the Lesser GNU General Public License as published
// by the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// This source file is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <http://www.gnu.org/licenses/>.
//
//
/////////////////////////////////////////////////////////////////////////

module floppy_track
(
	input         clk,
	input         reset,

	output [31:0] sd_lba,
	output reg    sd_rd,
	output reg    sd_wr,
	input         sd_ack,

	input   [8:0] sd_buff_addr,
	input   [7:0] sd_buff_dout,
	output  [7:0] sd_buff_din,
	input         sd_buff_wr,

	input         change,
	input         mount,
	input   [5:0] track,
	output reg    ready = 0,
	input         active,

	input  [12:0] ram_addr,
	output  [7:0] ram_do,
	input   [7:0] ram_di,
	input         ram_we,
	output reg    busy
);

assign sd_lba = lba;

reg  [31:0] lba;
reg   [3:0] rel_lba;

always @(posedge clk) begin
	reg old_ack;
	reg [5:0] cur_track ;
	reg old_change;
	reg saving ;
	reg dirty ;

	old_change <= change;
	old_ack <= sd_ack;

    if(sd_ack) {sd_rd,sd_wr} <= 0;

    if(ready && ram_we) dirty <= 1;
`ifdef SIMULATION
    if (sd_buff_wr & sd_ack) begin
        $display("FLOPPY DMA: write rel_lba=%0d addr=%03h data=%02h", rel_lba, sd_buff_addr, sd_buff_dout);
    end
`endif
`ifdef SIMULATION
    if (change && ~old_change) begin
        $display("FLOPPY: change edge detected (mount=%0d)", mount);
    end
`endif

    if(~old_change & change) begin
        ready <= mount;
        cur_track <= 'b111111;
        busy  <= 0;
        sd_rd <= 0;
        sd_wr <= 0;
        saving<= 0;
        dirty <= 0;
`ifdef SIMULATION
        $display("FLOPPY: change-> ready=%0d", mount);
`endif
    end
	else
	if(reset) begin
		cur_track <= 'b111111;
		busy  <= 0;
		sd_rd <= 0;
		sd_wr <= 0;
		saving<= 0;
		dirty <= 0;
	end
	else

    if(busy) begin
        if(old_ack && ~sd_ack) begin
            if(rel_lba != 4'd12) begin
                lba <= lba + 1'd1;
                rel_lba <= rel_lba + 1'd1;
                if(saving) sd_wr <= 1;
                    else sd_rd <= 1;
            end
            else
            if(saving && (cur_track != track)) begin
                saving <= 0;
                cur_track <= track;
                rel_lba <= 0;
                lba <= track * 8'd13; //track size = 1a00h = 13*512
                sd_rd <= 1;
            end
            else
            begin
                busy <= 0;
                dirty <= 0;
            end
        end
    end
    else
    // Only reload track when:
    // 1. Track changed AND drive is NOT active (don't interrupt reads/writes)
    // 2. Disk changed
    // 3. Dirty and inactive (save data)
    if(ready && (((cur_track != track) && ~active) || (old_change && ~change) || (dirty && ~active)))
        if (dirty && cur_track != 'b111111) begin
            saving <= 1;
            lba <= cur_track * 8'd13;
            rel_lba <= 0;
            sd_wr <= 1;
            busy <= 1;
        end
        else
        begin
            saving <= 0;
            cur_track <= track;
            rel_lba <= 0;
            lba <= track * 8'd13; //track size = 1a00h
            sd_rd <= 1;
            busy <= 1;
            dirty <= 0;
`ifdef SIMULATION
            $display("FLOPPY: load track %0d (LBA base=%0d) cur_track=%0d track_diff=%0d dirty=%0d active=%0d [track_input=%b]",
                     track, track*13, cur_track, (cur_track != track), dirty, active, track);
`endif
        end
end

/*
dpram #(13,8) floppy_dpram
(
        .clock_a(clk),
        .address_a({rel_lba, sd_buff_addr}),
        .wren_a(sd_buff_wr & sd_ack),
        .data_a(sd_buff_dout),
        .q_a(sd_buff_din),

        .clock_b(clk),
        .address_b(ram_addr),
        .wren_b(ram_we),
        .data_b(ram_di),
        .q_b(ram_do)

);
*/

bram #(.width_a(8),.widthad_a(13)) floppy_dpram 
(
        .clock_a(clk),
        .address_a({rel_lba, sd_buff_addr}),
        .wren_a(sd_buff_wr & sd_ack),
        .data_a(sd_buff_dout),
        .q_a(sd_buff_din),
        //.byteena_a(1'b1),

        .clock_b(clk),
        .address_b(ram_addr),
        .wren_b(ram_we),
        .data_b(ram_di),
        .q_b(ram_do),
        //.byteena_b(1'b1),
        .enable_a(1'b1),
        .enable_b(1'b1)
);

`ifdef SIMULATION
reg [12:0] prev_ram_addr;
reg prev_ram_we;
always @(posedge clk) begin
    prev_ram_addr <= ram_addr;
    prev_ram_we <= ram_we;
    // Debug track memory reads
    if (ram_addr != prev_ram_addr && !ram_we) begin
        $display("FTRACK: READ addr=%04h -> %02h", ram_addr, ram_do);
    end
    // Debug track memory writes
    if (ram_we && !prev_ram_we) begin
        $display("FTRACK: WRITE addr=%04h <- %02h", ram_addr, ram_di);
    end
end
`endif


/*
// Dual port track buffer
reg   [7:0] track_ram[13*512];

// IO controller side
always @(posedge clk) begin
	sd_buff_din <= track_ram[{rel_lba, sd_buff_addr}];
	if (sd_buff_wr & sd_ack) track_ram[{rel_lba, sd_buff_addr}] <= sd_buff_dout;
end

// Disk controller side
always @(posedge clk) begin
	ram_do <= track_ram[ram_addr];
	if (ram_we) track_ram[ram_addr] <= ram_di;
end
*/
endmodule
