import P65C816_pkg::*;

module mcode
  (
   input       CLK,
   input       RST_N,
   input       EN,
   input [7:0] IR,
   input [3:0] STATE,
   output MCode_r   M
   );
localparam logic [52:0] M_TAB[0:2047] = '{
// 00 BRK
{3'b111, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['PC++']
{3'b000, 4'b1100, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b100, 2'b10}, // ['PBR->[00:SP--]']
{3'b000, 4'b1100, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b010, 2'b10}, // ['PCH->[00:SP--]']
{3'b000, 4'b1100, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b010, 2'b10}, // ['PCL->[00:SP--]']
{3'b000, 4'b1100, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b001, 2'b10}, // ['P->[00:SP--]']
{3'b000, 4'b1111, 2'b00, 3'b010, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b10, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['[00:VECT+0]->DR', '00->PBR', '1->I']
{3'b010, 4'b1111, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b010, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10}, // ['[00:VECT+1]:DR->PC']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 01 ORA (DP,X)
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DX+X->DX']
{3'b000, 4'b0111, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[DX+0]->AAL']
{3'b000, 4'b0111, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[DX+1]->AAH']
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10}, // ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10}, // ['ALU([DBR:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 02 COP
{3'b111, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['PC++']
{3'b000, 4'b1000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b100, 2'b10}, // ['PBR->[00:SP--]']
{3'b000, 4'b1000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b010, 2'b10}, // ['PCH->[00:SP--]']
{3'b000, 4'b1000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b010, 2'b10}, // ['PCL->[00:SP--]']
{3'b000, 4'b1000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b001, 2'b10}, // ['P->[00:SP--]']
{3'b000, 4'b1111, 2'b00, 3'b010, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b10, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['[00:VECT+0]->DR', '00->PBR', '1->I']
{3'b010, 4'b1111, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b010, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10}, // ['[00:VECT+1]:DR->PC']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 03 ORA S
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['SPL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['SPH+Carry->DH']
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10}, // ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10}, // ['ALU([00:DX+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 04 TSB DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b110, 4'b0011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['[00:DX+0]->TL']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10}, // ['[00:DX+1]->TH']
{3'b110, 4'b0011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01111, 2'b11, 3'b000, 2'b00}, // ['ALU(T)->T', 'Flags']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10}, // ['TH->[00:DX+1]']
{3'b010, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['TL->[00:DX+0]']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 05 ORA DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10}, // ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10}, // ['ALU([00:DX+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 06 ASL DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b110, 4'b0011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['[00:DX+0]->TL']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10}, // ['[00:DX+1]->TH']
{3'b110, 4'b0011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01010, 2'b11, 3'b000, 2'b00}, // ['ALU(T)->T', 'Flags']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10}, // ['TH->[00:DX+1]']
{3'b010, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['TL->[00:DX+0]']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 07 ORA [DP]
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+0]->AAL']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+1]->AAH']
{3'b000, 4'b0011, 2'b10, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+2]->AB']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 08 PHP
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // []
{3'b010, 4'b1100, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b001, 2'b10}, // ['P->[00:SP--]']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 09 ORA IMM
{3'b100, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b01}, // ['ALU([PBR:PC])->AL', '[PBR:PC]->DR', 'PC++', 'Flags']
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b01}, // ['ALU([PBR:PC]:DR)->A', 'PC++', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 0A ASL A
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000010, 5'b01010, 2'b11, 3'b000, 2'b00}, // ['ALU(A)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 0B PHD
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // []
{3'b000, 4'b1000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b011000, 5'b00000, 2'b10, 3'b101, 2'b10}, // ['DH->[00:SP]', 'SP--']
{3'b010, 4'b1000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b011000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['DL->[00:SP]', 'SP--']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 0C TSB ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++']
{3'b110, 4'b0001, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['[DBR:AA+0]->TL']
{3'b000, 4'b0001, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10}, // ['[DBR:AA+1]->TH']
{3'b110, 4'b0001, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01111, 2'b11, 3'b000, 2'b00}, // ['ALU(T)->T', 'Flags']
{3'b000, 4'b0001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10}, // ['TH->[DBR:AA+1]']
{3'b010, 4'b0001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['TL->[DBR:AA+0]']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 0D ORA ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++']
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10}, // ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10}, // ['ALU([DBR:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 0E ASL ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++']
{3'b110, 4'b0001, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['[DBR:AA+0]->TL']
{3'b000, 4'b0001, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10}, // ['[DBR:AA+1]->TH']
{3'b110, 4'b0001, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01010, 2'b11, 3'b000, 2'b00}, // ['ALU(T)->T', 'Flags']
{3'b000, 4'b0001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10}, // ['TH->[DBR:AA+1]']
{3'b010, 4'b0001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['TL->[DBR:AA+0]']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 0F ORA LONG
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AB', 'PC++']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 10 BPL
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->DR', 'PC++']
{3'b011, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b100, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['PC+DR->PC']
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // []
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 11 ORA (DP), Y
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+0]->AAL', 'DBR->AB']
{3'b001, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+1]->AAH','AAL+YL->AAL']
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['AAH+YH+AALCarry->AAH']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 12 ORA (DP)
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+0]->AAL']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+1]->AAH']
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10}, // ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10}, // ['ALU([DBR:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 13 ORA (S),Y
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['SPL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['SPH+Carry->DH']
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+0]->AAL', 'DBR->AB']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+1]->AAH', 'AAL+YL->AAL']
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['AAH+YH+AALCarry->AAH']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 14 TRB DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b110, 4'b0011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['[00:DX+0]->TL']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10}, // ['[00:DX+1]->TH']
{3'b110, 4'b0011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01110, 2'b11, 3'b000, 2'b00}, // ['ALU(T)->T', 'Flags']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10}, // ['TH->[00:DX+1]']
{3'b010, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['TL->[00:DX+0]']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 15 ORA DP,X
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DX+Carry->DX']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DX+X->DX']
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10}, // ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10}, // ['ALU([00:DX+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 16 ASL DP,X
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DX+X->DX']
{3'b110, 4'b0011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['[00:DX+0]->TL']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10}, // ['[00:DX+1]->TH']
{3'b110, 4'b0011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01010, 2'b11, 3'b000, 2'b00}, // ['ALU(T)->T', 'Flags']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10}, // ['TH->[00:DX+1]']
{3'b010, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['TL->[00:DX+0]']
// 17 ORA [DP],Y
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+0]->AAL']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+1]->AAH','AAL+YL->AAL']
{3'b000, 4'b0011, 2'b10, 3'b000, 2'b00, 2'b01, 8'b00000101, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+2]->AB','AAH+YH+AALCarry->AAH']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 18 CLC
{3'b010, 4'b0000, 2'b00, 3'b100, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 19 ORA ABS,Y
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'DBR->AB', 'PC++']
{3'b001, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'AAL+XL/YL->AAL', 'PC++']
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['AAH+XH/YH+AALCarry->AAH']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 1A INC A
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000010, 5'b00011, 2'b11, 3'b000, 2'b00}, // ['ALU(A)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 1B TCS
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b100, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['A->S']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 1C TRB ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++']
{3'b110, 4'b0001, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['[DBR:AA+0]->TL']
{3'b000, 4'b0001, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10}, // ['[DBR:AA+1]->TH']
{3'b110, 4'b0001, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01110, 2'b11, 3'b000, 2'b00}, // ['ALU(T)->T', 'Flags']
{3'b000, 4'b0001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10}, // ['TH->[DBR:AA+1]']
{3'b010, 4'b0001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['TL->[DBR:AA+0]']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 1D ORA ABS,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'DBR->AB', 'PC++']
{3'b001, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'AAL+XL/YL->AAL', 'PC++']
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['AAH+XH/YH+AALCarry->AAH']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 1E ASL ABS,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'DBR->AB', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'AAL+XL/YL->AAL', 'PC++']
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['AAH+XH/YH+AALCarry->AAH']
{3'b110, 4'b0101, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['[AB:AA+0]->TL']
{3'b000, 4'b0101, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10}, // ['[AB:AA+1]->TH']
{3'b110, 4'b0101, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01010, 2'b11, 3'b000, 2'b00}, // ['ALU(T)->T', 'Flags']
{3'b000, 4'b0101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10}, // ['TH->[AB:AA+1]']
{3'b010, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['TL->[AB:AA+0]']
// 1F ORA LONG,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'AAL+XL/YL->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000101, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AB', 'AAH+XH/YH+AALCarry->AAH', 'PC++']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 20 JSR ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL, 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // []
{3'b000, 4'b1100, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b010, 2'b10}, // ['PCH->[00:SP]', 'SP--']
{3'b010, 4'b1100, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b110, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b010, 2'b10}, // ['PCL->[00:SP]', 'SP--', 'AA->PC']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 21 AND (DP,X)
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DX+X->DX']
{3'b000, 4'b0111, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+0]->AAL']
{3'b000, 4'b0111, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+1]->AAH']
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10}, // ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10}, // ['ALU([DBR:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 22 JSR LONG
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++']
{3'b000, 4'b1000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b100, 2'b10}, // ['PBR->[00:SP]', 'SP--']
{3'b000, 4'b1000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // []
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b10, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->PBR']
{3'b000, 4'b1000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b010, 2'b10}, // ['PCH->[00:SP]', 'SP--']
{3'b010, 4'b1000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b110, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b010, 2'b10}, // ['PCL->[00:SP]', 'SP--', 'AA->PC']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 23 AND S
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['SPL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['SPH+Carry->DH']
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10}, // ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10}, // ['ALU([00:DX+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 24 BIT DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b01001, 2'b01, 3'b000, 2'b10}, // ['ALU([00:DX+0])', '[00:DX+0]->DR', 'Flags']
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b01001, 2'b10, 3'b000, 2'b10}, // ['ALU([00:DX+1]:DR)', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 25 AND DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10}, // ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10}, // ['ALU([00:DX+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 26 ROL DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b110, 4'b0011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['[00:DX+0]->TL']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10}, // ['[00:DX+1]->TH']
{3'b110, 4'b0011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01100, 2'b11, 3'b000, 2'b00}, // ['ALU(T)->T', 'Flags']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10}, // ['TH->[00:DX+1]']
{3'b010, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['TL->[00:DX+0]']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 27 AND [DP]
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+0]->AAL']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+1]->AAH']
{3'b000, 4'b0011, 2'b10, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+2]->AB']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 28 PLP
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // []
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['SP++']
{3'b010, 4'b1100, 2'b00, 3'b011, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[SP]->P', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 29 AND IMM
{3'b100, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b01}, // ['ALU([PBR:PC])->AL', '[PBR:PC]->DR', 'PC++', 'Flags']
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b01}, // ['ALU([PBR:PC]:DR)->A', 'PC++', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 2A ROL A
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000010, 5'b01100, 2'b11, 3'b000, 2'b00}, // ['ALU(A)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 2B PLD
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // []
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b110, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['SP++']
{3'b000, 4'b1000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b110, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['[00:SP++]->DR']
{3'b010, 4'b1000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b01, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10}, // ['ALU([00:SP]:DR)->D', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 2C BIT ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++']
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b01001, 2'b01, 3'b000, 2'b10}, // ['ALU([DBR:AA+0])', '[DBR:AA+0]->DR', 'Flags']
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b01001, 2'b10, 3'b000, 2'b10}, // ['ALU([DBR:AA+1]:DR)', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 2D AND ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++']
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10}, // ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10}, // ['ALU([DBR:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 2E ROL ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++']
{3'b110, 4'b0001, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['[DBR:AA+0]->TL']
{3'b000, 4'b0001, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10}, // ['[DBR:AA+1]->TH']
{3'b110, 4'b0001, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01100, 2'b11, 3'b000, 2'b00}, // ['ALU(T)->T', 'Flags']
{3'b000, 4'b0001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10}, // ['TH->[DBR:AA+1]']
{3'b010, 4'b0001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['TL->[DBR:AA+0]']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 2F AND LONG
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AB', 'PC++']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A, 'Flags'']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 30 BMI
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->DR', 'PC++']
{3'b011, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b100, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['PC+DR->PC']
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // []
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 31 AND (DP),Y
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+0]->AAL', 'DBR->AB']
{3'b001, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+1]->AAH', 'AAL+YL->AAL ']
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['AAH+YH+AALCarry->AAH']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 32 AND (DP)
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+0]->AAL']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+1]->AAH']
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10}, // ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10}, // ['ALU([DBR:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 33 AND (S),Y
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['SPL+[PBR:PC]->DX', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+0]->AAL', 'DBR->AB']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+1]->AAH', 'AAL+Y->AAL']
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['AAH+YH+AALCarry->AAH']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 34 BIT DP,X
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DX+Carry->DX']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DX+X->DX']
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b01001, 2'b01, 3'b000, 2'b10}, // ['ALU([00:DX+0]', '[00:DX+0]->DR', 'Flags']
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b01001, 2'b10, 3'b000, 2'b10}, // ['ALU([00:DX+1]', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 35 AND DP,X
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DX+Carry->DX']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DX+X->DX']
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10}, // ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10}, // ['ALU([00:DX+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 36 ROL DP,X
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DX+X->DX']
{3'b110, 4'b0011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['[00:DX+0]->TL']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10}, // ['[00:DX+1]->TH']
{3'b110, 4'b0011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01100, 2'b11, 3'b000, 2'b00}, // ['ALU(T)->T', 'Flags']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10}, // ['TH->[00:DX+1]']
{3'b010, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['TL->[00:DX+0]']
// 37 AND [DP],Y
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+0]->AAL']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+1]->AAH,AAL+Y->AAL']
{3'b000, 4'b0011, 2'b10, 3'b000, 2'b00, 2'b01, 8'b00000101, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+2]->AB','AAH+YH+AALCarry->AAH']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 38 SEC
{3'b010, 4'b0000, 2'b00, 3'b100, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 39 AND ABS,Y
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'DBR->AB', 'PC++']
{3'b001, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'AAL+XL/YL->AAL', 'PC++']
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['AAH+XH/YH+AALCarry->AAH']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 3A DEC A
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000010, 5'b00010, 2'b11, 3'b000, 2'b00}, // ['ALU(A)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 3B TSC
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b101010, 5'b00001, 2'b11, 3'b000, 2'b00}, // ['ALU(SP)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 3C BIT ABS,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
{3'b001, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL']
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['AAH+XH/YH+AALCarry->AAH']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b01001, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b01001, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1])' 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 3D AND ABS,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'DBR->AB', 'PC++']
{3'b001, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'AAL+XL/YL->AAL', 'PC++']
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['AAH+XH/YH+AALCarry->AAH']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 3E ROL ABS, X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'DBR->AB', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'AAL+XL/YL->AAL', 'PC++']
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['AAH+XH/YH+AALCarry->AAH'']
{3'b110, 4'b0101, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['[AB:AA+0]->TL']
{3'b000, 4'b0101, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10}, // ['[AB:AA+1]->TH']
{3'b110, 4'b0101, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01100, 2'b11, 3'b000, 2'b00}, // ['ALU(T)->T', 'Flags']
{3'b000, 4'b0101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10}, // ['TH->[AB:AA+1]']
{3'b010, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['TL->[AB:AA+0]']
// 3F AND LONG,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'AAL+XL/YL->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000101, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AB', 'AAH+XH/YH+AALCarry->AAH', 'PC++']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 40 RTI
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['SP++']
{3'b000, 4'b1100, 2'b00, 3'b011, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:SP]->P', 'SP++']
{3'b000, 4'b1100, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:SP]->DR', 'SP++']
{3'b111, 4'b1100, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b010, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:SP]:DR->PC']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['SP++']
{3'b010, 4'b1100, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b10, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:SP]->PBR']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 41 EOR (DP,X)
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DX+X->DX']
{3'b000, 4'b0111, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+0]->AAL']
{3'b000, 4'b0111, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+1]->AAH']
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10}, // ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10}, // ['ALU([DBR:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 42 WDM
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['PC++']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 43 EOR S
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['SPL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10}, // ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10}, // ['ALU([00:DX+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 44 MVP
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b11, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->DBR', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b10, 8'b00000001, 3'b001, 3'b000, 3'b110, 2'b00, 6'b001010, 5'b00010, 2'b11, 3'b000, 2'b01}, // ['[PBR:PC]->ABR', 'PC++', 'X->AA', 'X-1->X']
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b11, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b010010, 5'b00010, 2'b11, 3'b000, 2'b10}, // ['[ABR:AA]->DR', 'Y->AA', 'Y-1->Y']
{3'b000, 4'b0001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b110, 2'b10}, // ['DR->[DBR:AA]']
{3'b000, 4'b0001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b111, 3'b000, 3'b101, 2'b00, 6'b000101, 5'b10000, 2'b11, 3'b000, 2'b00}, // ['ALU(A)->A', 'PC-3->PC']
{3'b010, 4'b0001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // []
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 45 EOR DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10}, // ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10}, // ['ALU([00:DX+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 46 LSR DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b110, 4'b0011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['[00:DX+0]->TL']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10}, // ['[00:DX+1]->TH']
{3'b110, 4'b0011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01011, 2'b11, 3'b000, 2'b00}, // ['ALU(T)->T', 'Flags']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10}, // ['TH->[00:DX+1]']
{3'b010, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['TL->[00:DX+0]']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 47 EOR [DP]
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+0]->AAL']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+1]->AAH']
{3'b000, 4'b0011, 2'b10, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+2]->AB']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 48 PHA
{3'b110, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // []
{3'b000, 4'b1100, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b001, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b101, 2'b10}, // ['AH->[00:SP]', 'SP--']
{3'b010, 4'b1100, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b001, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['AL->[00:SP]', 'SP--']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 49 EOR IMM
{3'b100, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b01}, // ['ALU([PBR:PC])->AL', '[PBR:PC]->DR', 'PC++', 'Flags']
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b01}, // ['ALU([PBR:PC]:DR)->A', 'PC++', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 4A LSR A
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000010, 5'b01011, 2'b11, 3'b000, 2'b00}, // ['ALU(REG+1)->REG', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 4B PHK
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // []
{3'b010, 4'b1100, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b110000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['PBR->[00:SP]', 'SP--']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 4C JMP ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->DR', 'PC++']
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b010, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]:DR->PC']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 4D EOR ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++']
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10}, // ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10}, // ['ALU([DBR:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 4E LSR ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++']
{3'b110, 4'b0001, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['[DBR:AA+0]->TL']
{3'b000, 4'b0001, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10}, // ['[DBR:AA+1]->TH']
{3'b110, 4'b0001, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01011, 2'b11, 3'b000, 2'b00}, // ['ALU(T)->T', 'Flags']
{3'b000, 4'b0001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10}, // ['TH->[DBR:AA+1]']
{3'b010, 4'b0001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['TL->[DBR:AA+0]']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 4F EOR LONG
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AB', 'PC++']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 50 BVC
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->DL', 'PC++']
{3'b011, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b100, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['PC+DL->PC']
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['NOP']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 51 EOR (DP),Y
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+0]->AAL', 'DBR->AB']
{3'b001, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+1]->AAH', 'AAL+YL->AAL ']
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['AAH+YH+AALCarry->AAH']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 52 EOR (DP)
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // [00:DX+0]->AAL
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // [00:DX+1]->AAH
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10}, // ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10}, // ['ALU([DBR:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 53 EOR (S),Y
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['SPL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+0]->AAL', 'DBR->AB']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+1]->AAH', 'AAL+YL->AAL ']
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['AAH+YH+AALCarry->AAH']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 54 MVN
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b11, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->DBR', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b10, 8'b00000001, 3'b001, 3'b000, 3'b110, 2'b00, 6'b001010, 5'b00011, 2'b11, 3'b000, 2'b01}, // ['[PBR:PC]->ABR', 'PC++', 'X->AA', 'X+1->X']
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b11, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b010010, 5'b00011, 2'b11, 3'b000, 2'b10}, // ['[ABR:AA]->DR', 'Y->AA', 'Y+1->Y']
{3'b000, 4'b0001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b110, 2'b10}, // ['DR->[DBR:AA]']
{3'b000, 4'b0001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b111, 3'b000, 3'b101, 2'b00, 6'b000101, 5'b10000, 2'b11, 3'b000, 2'b00}, // ['ALU(A-1)->A','PC-3->PC']
{3'b010, 4'b0001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // []
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 55 EOR DP,X
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DX+Carry->DX']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DX+X->DX']
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10}, // ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10}, // ['ALU([00:DX+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 56 LSR DP,X
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DX+X->DX']
{3'b110, 4'b0011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['[00:DX+0]->TL']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10}, // ['[00:DX+1]->TH']
{3'b110, 4'b0011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01011, 2'b11, 3'b000, 2'b00}, // ['ALU(T)->T', 'Flags']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10}, // ['TH->[00:DX+1]']
{3'b010, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['TL->[00:DX+0]']
// 57 EOR [DP],Y
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+0]->AAL']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+1]->AAH,AAL+YL->AAL']
{3'b000, 4'b0011, 2'b10, 3'b000, 2'b00, 2'b01, 8'b00000101, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+2]->AB','AAH+YH+AALCarry->AAH']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 58 CLI
{3'b010, 4'b0000, 2'b00, 3'b100, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['[PBR:PC]->,ALU()->A', 'Flags', 'ALU()->X,Y', 'ALU()->A']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 59 EOR ABS,Y
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
{3'b001, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL']
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['AAH+XH/YH+AALCarry->AAH']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 5A PHY
{3'b110, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b011, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // []
{3'b000, 4'b1100, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b011, 2'b00, 6'b010000, 5'b00000, 2'b10, 3'b101, 2'b10}, // ['YH->[00:SP]', 'SP--']
{3'b010, 4'b1100, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b011, 2'b00, 6'b010000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['YL->[00:SP]', 'SP--']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 5B TCD
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b01, 6'b000010, 5'b00001, 2'b00, 3'b000, 2'b00}, // ['ALU(A)->D', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 5C JMP LONG
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++']
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b110, 3'b000, 3'b000, 2'b10, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->PBR', 'AA->PC']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 5D EOR ABS,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
{3'b001, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL']
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['AAH+XH/YH+AALCarry->AAH']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 5E LSR ABS,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL']
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['AAH+XH/YH+AALCarry->AAH']
{3'b110, 4'b0101, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['[AB:AA+0]->TL']
{3'b000, 4'b0101, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10}, // ['[AB:AA+1]->TH']
{3'b110, 4'b0101, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01011, 2'b11, 3'b000, 2'b00}, // ['ALU(T)->T', 'Flags']
{3'b000, 4'b0101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10}, // ['TH->[AB:AA+1]']
{3'b010, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['TL->[AB:AA+0]']
// 5F EOR LONG,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000101, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AB', 'PC++', 'AAH+XH/YH+AALCarry->AAH']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 60 RTS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['SP++']
{3'b000, 4'b1100, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:SP]->DR', 'SP++']
{3'b000, 4'b1100, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b010, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:SP]:DR->PC']
{3'b010, 4'b1100, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['PC++']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 61 ADC (DP,X)
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DX+X->DX']
{3'b000, 4'b0111, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+0]->AAL']
{3'b000, 4'b0111, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+1]->AAH']
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10}, // ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10}, // ['ALU([DBR:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 62 PER
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->TL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->TH', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01101100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['PC+Offset->AA']
{3'b000, 4'b1000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b011, 2'b10}, // ['AAH->[00:SP]', 'SP--']
{3'b010, 4'b1000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b011, 2'b10}, // ['AAL->[00:SP]', 'SP--']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 63 ADC S
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['SPL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10}, // ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10}, // ['ALU([00:DX+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 64 STZ DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b100, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b111, 2'b10}, // ['0->[00:DX+0]']
{3'b010, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b111, 2'b10}, // ['0->[00:DX+1]']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 65 ADC DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10}, // ['[00:DX+0]->A']
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10}, // ['[00:DX+1]->A']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 66 ROR DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b110, 4'b0011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['[00:DX+0]->TL']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10}, // ['[00:DX+1]->TH']
{3'b110, 4'b0011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01101, 2'b11, 3'b000, 2'b00}, // ['ALU(T)->T', 'Flags']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10}, // ['TH->[00:DX+1]']
{3'b010, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['TL->[00:DX+0]']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 67 ADC [DP]
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+0]->AAL']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+1]->AAH']
{3'b000, 4'b0011, 2'b10, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+2]->AB']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 68 PLA
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, //
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['SP++']
{3'b100, 4'b1100, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b010, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['ALU([00:SP])->REGL', 'SP++']
{3'b010, 4'b1100, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10}, // ['ALU([00:SP])->REGH']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 69 ADC IMM
{3'b100, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b01}, // ['ALU([PBR:PC])->AL', '[PBR:PC]->DR', 'PC++', 'Flags']
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b01}, // ['ALU([PBR:PC]:DR)->A', 'PC++', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 6A ROR A
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000010, 5'b01101, 2'b11, 3'b000, 2'b00}, // ['ALU(REG+1)->REG', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 6B RTL
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['SP++']
{3'b000, 4'b1000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:SP]->DR', 'SP++']
{3'b000, 4'b1000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b010, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:SP]:DR->PC', 'SP++']
{3'b010, 4'b1000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b10, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:SP]->PBR', 'PC++']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 6C JMP (ABS)
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++']
{3'b000, 4'b0110, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:AA+0]->DR']
{3'b010, 4'b0110, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b010, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:AA+1]:DR->PC']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 6D ADC ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++']
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10}, // ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10}, // ['ALU([DBR:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 6E ROR ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++']
{3'b110, 4'b0001, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['[DBR:AA+0]->TL']
{3'b000, 4'b0001, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10}, // ['[DBR:AA+1]->TH']
{3'b110, 4'b0001, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01101, 2'b11, 3'b000, 2'b00}, // ['ALU(T)->T', 'Flags']
{3'b000, 4'b0001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10}, // ['TH->[DBR:AA+1]']
{3'b010, 4'b0001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['TL->[DBR:AA+0]']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 6F ADC LONG
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AB', 'PC++']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 70 BVS
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->DR', 'PC++']
{3'b011, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b100, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['PC+DR->PC']
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // []
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 71 ADC (DP),Y
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+0]->AAL', 'DBR->AB']
{3'b001, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+1]->AAH', 'AAL+YL->AAL ']
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['AAH+YH+AALCarry->AAH']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 72 ADC (DP)
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // [00:DX+0]->AAL
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // [00:DX+1]->AAH
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10}, // ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10}, // ['ALU([DBR:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 73 ADC (S),Y
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['SPL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+0]->AAL', 'DBR->AB']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+1]->AAH', 'AAL+YL->AAL']
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['AAH+YH+AALCarry->AAH']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 74 STZ DP,X
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DX+X->DX']
{3'b100, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b111, 2'b10}, // ['0->[00:DX+0]']
{3'b010, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b111, 2'b10}, // ['0->[00:DX+1]']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 75 ADC DP,X
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DX+Carry->DX']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DX+X->DX']
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10}, // ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10}, // ['ALU([00:DX+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 76 ROR DP,X
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DX+X->DX']
{3'b110, 4'b0011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['[00:DX+0]->TL']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10}, // ['[00:DX+1]->TH']
{3'b110, 4'b0011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01101, 2'b11, 3'b000, 2'b00}, // ['ALU(T)->T', 'Flags']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10}, // ['TH->[00:DX+1]']
{3'b010, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10}, // ['TL->[00:DX+0]']
// 77 ADC [DP],Y
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+0]->AAL']
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+1]->AAH', 'AAL+YL->AAL']
{3'b000, 4'b0011, 2'b10, 3'b000, 2'b00, 2'b01, 8'b00000101, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10}, // ['[00:DX+2]->AB', 'AAH+YH+AALCarry->AAH']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 78 SEI
{3'b010, 4'b0000, 2'b00, 3'b100, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['[PBR:PC]->,ALU()->A', 'Flags', 'ALU()->X,Y', 'ALU()->A']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 79 ADC ABS,Y
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
{3'b001, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL']
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['AAH+XH/YH+AALCarry->AAH']
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10}, // ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10}, // ['ALU([AB:AA+1]:DR)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 7A PLY
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // []
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['SP++']
{3'b100, 4'b1100, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b010, 3'b111, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10}, // ['ALU([00:SP])->YL', 'SP++']
{3'b010, 4'b1100, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10}, // ['ALU([00:SP])->YH']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 7B TDC
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b011010, 5'b00001, 2'b11, 3'b000, 2'b00}, // ['ALU(D)->A', 'Flags']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 7C JMP (ABS,X)
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['AAH+XH/YH+Carry->AAH']
{3'b000, 4'b0010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:AA+0]->DR']
{3'b010, 4'b0010, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b010, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:AA+1]:DR->PC']
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 7D ADC ABS,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 7E ROR ABS,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 4'b0101, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 4'b0101, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 4'b0101, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01101, 2'b11, 3'b000, 2'b00},
{3'b000, 4'b0101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
// 7F ADC LONG,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000101, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 80 BRA
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['[PBR:PC]->DL', 'PC++']
{3'b011, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b100, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['PC+DL->PC']
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // []
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 81 STA (DP,X)
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0111, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0111, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 4'b0001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 4'b0001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 82 BRL
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01101100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b011, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 83 STA S
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 84 STY DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b011, 2'b00, 6'b010010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b011, 2'b00, 6'b010010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 85 STA DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01}, // ['DL+[PBR:PC]->DL', 'PC++']
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00}, // ['DH+Carry->DH']
{3'b100, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10}, // REGL->[00:DX+0]
{3'b010, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10}, // REGH->[D00:X+1]
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 86 STX DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b010, 2'b00, 6'b001010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b010, 2'b00, 6'b001010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 87 STA [DP]
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b10, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 88 DEY
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b010010, 5'b00010, 2'b11, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 89 BIT IMM
{3'b100, 4'b0000, 2'b00, 3'b111, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b01001, 2'b01, 3'b000, 2'b01},
{3'b010, 4'b0000, 2'b00, 3'b111, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b01001, 2'b10, 3'b000, 2'b01},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 8A TXA
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b001010, 5'b00000, 2'b11, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 8B PHB
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 4'b1100, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b111010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 8C STY ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 4'b0001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b011, 2'b00, 6'b010010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 4'b0001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b011, 2'b00, 6'b010010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 8D STA ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 4'b0001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 4'b0001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 8E STX ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 4'b0001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b010, 2'b00, 6'b001010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 4'b0001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b010, 2'b00, 6'b001010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 8F STA LONG
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 90 BCC
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b011, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b100, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 91 STA (DP),Y
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 92 STA (DP)
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 4'b0001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00100, 2'b01, 3'b101, 2'b10},
{3'b010, 4'b0001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 93 STA (S),Y
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 94 STY DP,X
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b011, 2'b00, 6'b010010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b011, 2'b00, 6'b010010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 95 STA DP,X
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 96 STX DP,Y
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b01, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b010, 2'b00, 6'b001010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b010, 2'b00, 6'b001010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 97 STA [DP],Y
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b10, 3'b000, 2'b00, 2'b01, 8'b00000101, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 98 TYA
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b010010, 5'b00000, 2'b11, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 99 STA ABS,Y
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 9A TXS
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b101, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 9B TXY
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b001010, 5'b00000, 2'b11, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 9C STZ ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 4'b0001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b111, 2'b10},
{3'b010, 4'b0001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b111, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 9D STA ABS,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 9E STZ ABS,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b111, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b111, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// 9F STA LONG,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000101, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// A0 LDY IMM
{3'b100, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b111, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b01},
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b111, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b01},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// A1 LDA (DP,X)
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0111, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0111, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// A2 LDX IMM
{3'b100, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b110, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b01},
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b110, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b01},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// A3 LDA S
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// A4 LDY DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// A5 LDA DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// A6 LDX DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// A7 LDA [DP]
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b10, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// A8 TAY
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b000010, 5'b00000, 2'b11, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// A9 LDA IMM
{3'b100, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b01},
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b01},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// AA TAX
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b000010, 5'b00000, 2'b11, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// AB PLB
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 4'b1000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b11, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// AC LDY ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// AD LDA ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// AE LDX ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// AF LDA LONG
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// B0 BCS
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b011, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b100, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// B1 LDA (DP),Y
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b001, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// B2 LDA (DP)
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// B3 LDA (S),Y
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// B4 LDY DP,X
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// B5 LDA DP,X
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// B6 LDX DP,Y
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b01, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// B7 LDA [DP],Y
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b10, 3'b000, 2'b00, 2'b01, 8'b00000101, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// B8 CLV
{3'b010, 4'b0000, 2'b00, 3'b100, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// B9 LDA ABS,Y
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// BA TSX
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b101010, 5'b00001, 2'b11, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// BB TYX
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b010010, 5'b00000, 2'b11, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// BC LDY ABS,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// BD LDA ABS,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// BE LDX ABS,Y
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// BF LDA LONG,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000101, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// C0 CPY IMM
{3'b100, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b011, 2'b00, 6'b010000, 5'b10000, 2'b01, 3'b000, 2'b01},
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b011, 2'b00, 6'b010001, 5'b10000, 2'b10, 3'b000, 2'b01},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// C1 CMP (DP,X)
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0111, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0111, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// C2 REP
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b010, 4'b0000, 2'b00, 3'b110, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// C3 CMP S
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// C4 CPY DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b011, 2'b00, 6'b010000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b011, 2'b00, 6'b010001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// C5 CMP DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// C6 DEC DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 4'b0011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 4'b0011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100010, 5'b00010, 2'b11, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// C7 CMP [DP]
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b10, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// C8 INY
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b010010, 5'b00011, 2'b11, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// C9 CMP IMM
{3'b100, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b01},
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b01},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// CA DEX
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b001010, 5'b00010, 2'b11, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// CB WAI
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// CC CPY ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b011, 2'b00, 6'b010000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b011, 2'b00, 6'b010001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// CD CMP ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// CE DEC ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b110, 4'b0001, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 4'b0001, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 4'b0001, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100010, 5'b00010, 2'b11, 3'b000, 2'b00},
{3'b000, 4'b0001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 4'b0001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// CF CMP LONG
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// D0 BNE
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b011, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b100, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// D1 CMP (DP),Y
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b001, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// D2 CMP (DP)
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// D3 CMP (S),Y
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// D4 PEI
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b1000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b011, 2'b10},
{3'b010, 4'b1000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b011, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// D5 CMP DP,X
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// D6 DEC DP,X
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 4'b0011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 4'b0011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100010, 5'b00010, 2'b11, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
// D7 CMP [DP],Y
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b10, 3'b000, 2'b00, 2'b01, 8'b00000101, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// D8 CLD
{3'b010, 4'b0000, 2'b00, 3'b100, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// D9 CMP ABS,Y
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// DA PHX
{3'b110, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b010, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b1100, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b010, 2'b00, 6'b001000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 4'b1100, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b010, 2'b00, 6'b001000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// DB STP
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// DC JMP [ABS]
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0110, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0110, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b010, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b010, 4'b0110, 2'b10, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b10, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// DD CMP ABS,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// DE DEC ABS,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 4'b0101, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 4'b0101, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 4'b0101, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100010, 5'b00010, 2'b11, 3'b000, 2'b00},
{3'b000, 4'b0101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
// DF CMP LONG,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000101, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// E0 CPX IMM
{3'b100, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b010, 2'b00, 6'b001000, 5'b10000, 2'b01, 3'b000, 2'b01},
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b010, 2'b00, 6'b001001, 5'b10000, 2'b10, 3'b000, 2'b01},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// E1 SBC (DP,X)
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0111, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0111, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// E2 SEP
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b010, 4'b0000, 2'b00, 3'b110, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// E3 SBC S
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// E4 CPX DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b010, 2'b00, 6'b001000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b010, 2'b00, 6'b001001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// E5 SBC DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// E6 INC DP
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 4'b0011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 4'b0011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100010, 5'b00011, 2'b11, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// E7 SBC [DP]
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b10, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// E8 INX
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b001010, 5'b00011, 2'b11, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// E9 SBC IMM
{3'b100, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b01},
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b01},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// EA NOP
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// EB XBA
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b11, 3'b000, 2'b00},
{3'b010, 4'b0000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// EC CPX ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b010, 2'b00, 6'b001000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b010, 2'b00, 6'b001001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// ED SBC ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// EE INC ABS
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b110, 4'b0001, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 4'b0001, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 4'b0001, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100010, 5'b00011, 2'b11, 3'b000, 2'b00},
{3'b000, 4'b0001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 4'b0001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// EF SBC LONG
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// F0 BEQ
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b011, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b100, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// F1 SBC (DP),Y
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b001, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// F2 SBC (DP)
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 4'b0001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// F3 SBC (S),Y
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// F4 PEA
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b1000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b011, 2'b10},
{3'b010, 4'b1000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b011, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// F5 SBC DP,X
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// F6 INC DP,X
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 4'b0011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 4'b0011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100010, 5'b00011, 2'b11, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
// F7 SBC [DP],Y
{3'b101, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 4'b0011, 2'b10, 3'b000, 2'b00, 2'b01, 8'b00000101, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// F8 SED
{3'b010, 4'b0000, 2'b00, 3'b100, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// F9 SBC ABS,Y
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// FA PLX
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b1100, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b010, 3'b110, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b1100, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// FB XCE
{3'b010, 4'b0000, 2'b00, 3'b101, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// FC JSR (ABS,X)
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b1000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b010, 2'b10},
{3'b000, 4'b1000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b010, 2'b10},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 4'b0010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b010, 4'b0010, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b010, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// FD SBC ABS,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
// FE INC ABS,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 4'b0101, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 4'b0101, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 4'b0101, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100010, 5'b00011, 2'b11, 3'b000, 2'b00},
{3'b000, 4'b0101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 4'b0101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
// FF SBC LONG,X
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000101, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 4'b0101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 4'b0101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 4'bXXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX}};

   localparam logic [7:0] ALU_TAB[0:16] = '{
      {3'b100, 3'b100, 1'b0, 1'b0},
      {3'b100, 3'b100, 1'b0, 1'b1},
      {3'b110, 3'b100, 1'b0, 1'b0},
      {3'b111, 3'b100, 1'b0, 1'b0},
      {3'b100, 3'b000, 1'b0, 1'b0},
      {3'b100, 3'b001, 1'b0, 1'b0},
      {3'b100, 3'b010, 1'b0, 1'b0},
      {3'b100, 3'b011, 1'b0, 1'b0},
      {3'b100, 3'b111, 1'b1, 1'b0},
      {3'b100, 3'b001, 1'b1, 1'b0},
      {3'b000, 3'b100, 1'b0, 1'b0},
      {3'b010, 3'b100, 1'b0, 1'b0},
      {3'b001, 3'b100, 1'b0, 1'b0},
      {3'b011, 3'b100, 1'b0, 1'b0},
      {3'b100, 3'b101, 1'b0, 1'b0},
      {3'b100, 3'b101, 1'b1, 1'b0},
      {3'b100, 3'b110, 1'b0, 1'b0}
   };

   MicroInst_r         MI;
   ALUCtrl_r        ALUFlags;

   assign ALUFlags = ALU_TAB[MI.ALUCtrl];


   always @(posedge CLK or negedge RST_N)
   begin: xhdl0
      reg [3:0]   STATE2;
      if (RST_N == 1'b0)
         MI <= {3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b11};
      else
      begin
         STATE2 = STATE - 1;
         if (EN == 1'b1)
         begin
            if (STATE == 4'b0000)
               MI <= {3'b000, 4'b0000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b11};
            else
              MI <= M_TAB[({IR, STATE2[2:0]})];
         end
      end
   end

   assign M = {ALUFlags, MI.stateCtrl, MI.addrBus, MI.addrInc, MI.muxCtrl, MI.addrCtrl, MI.loadPC, MI.loadSP, MI.regAXY, MI.loadP, MI.loadT, MI.loadDKB, MI.busCtrl, MI.byteSel, MI.outBus, MI.va};

endmodule
