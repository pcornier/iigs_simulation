//
// iwm_flux.v: IWM Core with Flux Transition Interface
//
// This module implements the IWM's flux decoding and register read logic.
// Soft switch state (Q6, Q7, phases, motor) is received as INPUTS from
// the parent module (iwm_woz.v), which is the single source of truth.
//
// Key responsibilities:
// - Flux transition decoding (window-based state machine)
// - Data/shift register management
// - Register read mux (data, status, handshake)
//
// Reference: MAME iwm.cpp (src/devices/machine/iwm.cpp)
//

// Enable detailed byte framing debug output for comparing with MAME
// Uncomment the following line to enable:
`define BYTE_FRAME_DEBUG

// Enable sector read logging with checksum validation
// Uncomment the following line to enable:
`define SECTOR_DEBUG

module iwm_flux (
    // Global signals
    input  wire        CLK_14M,         // 14MHz master clock
    input  wire        CLK_7M_EN,       // 7MHz clock enable (IWM runs at 7M like real hardware)
    input  wire        RESET,
    input  wire        CEN,             // Clock enable (phi2) for CPU bus timing

    // CPU interface
    input  wire [3:0]  ADDR,            // $C0E0-$C0EF offset (for register read mux)
    input  wire        RD,              // Read strobe (active high)
    input  wire        WR,              // Write strobe (active high)
    input  wire [7:0]  DATA_IN,         // Data from CPU (for mode register write)
    output wire [7:0]  DATA_OUT,        // Data to CPU

    // Soft switch state from iwm_woz.v (SINGLE SOURCE OF TRUTH)
    input  wire [3:0]  SW_PHASES,       // Current phase state
    input  wire        SW_MOTOR_ON,     // Motor on command
    input  wire        SW_DRIVE_SEL,    // Drive select
    input  wire        SW_Q6,           // Q6 latch state
    input  wire        SW_Q7,           // Q7 latch state
    input  wire [7:0]  SW_MODE,         // Mode register

    // Flux interface from drive (active high pulse when flux reversal detected)
    input  wire        FLUX_TRANSITION,

    // Status inputs from drive
    input  wire        MOTOR_ACTIVE,    // Motor command is on (like MAME m_active, not gated by disk)
    input  wire        MOTOR_SPINNING,  // Physical motor state (gated by disk presence, for byte decoding)
    input  wire        DISK_READY,      // Track data is valid and motor spinning
    input  wire        DISK_MOUNTED,    // Disk image is loaded (independent of motor)

    // Drive type selection
    input  wire        IS_35_INCH,      // 1 = 3.5" drive, 0 = 5.25" drive

    // Per-drive status sensing (computed by flux_drive, muxed by iwm_woz)
    input  wire        SENSE_BIT,       // Status sense from selected drive
    input  wire [2:0]  LATCHED_SENSE_REG, // Latched sense register index (for debug logging)
    input  wire        DISKREG_SEL,     // SEL bit from $C031 (for debug logging)

    // Disk position for debug logging (to compare with MAME)
    input  wire [16:0] DISK_BIT_POSITION, // Current bit position on track

    // Write output (future use)
    output wire        FLUX_WRITE,      // Pulse when writing flux transition

    // Debug
    output wire [7:0]  DEBUG_RSH,       // Read shift register (for debug)
    output wire [2:0]  DEBUG_STATE      // State machine state (for debug)
);

    //=========================================================================
    // IWM Data Registers
    //=========================================================================

    reg [7:0]  m_data;      // Data register - holds completed byte from disk
    reg [7:0]  m_rsh;       // Read shift register - bits shift in here
    reg [7:0]  m_wsh;       // Write shift register - bits shift out here
    reg [7:0]  m_whd;       // Write handshake register (MAME: initialized to 0xBF)
    reg        m_data_read; // Flag: data register has been read since last byte loaded
    reg        m_rw_mode;   // 0 = read mode, 1 = write mode (tracks Q7 for mode changes)
    reg        m_motor_was_on; // Track motor state for edge detection
    reg [5:0]  async_update;   // MAME: countdown to clear m_data in async mode (14 cycles at 7MHz = 2µs)
    reg        bit7_acknowledged; // MAME: bit 7 was read, mask it for subsequent reads
    reg        rd_latched;  // Edge detection: tracks if current RD has been processed

    // Async mode: mode bit 1 = 1 means async (MAME: is_sync() = !(mode & 0x02))
    wire       is_async = SW_MODE[1];

    //=========================================================================
    // State Machine (from MAME)
    //=========================================================================

    localparam S_IDLE           = 3'd0;
    localparam SR_WINDOW_EDGE_0 = 3'd1;  // Reading: waiting for flux transition
    localparam SR_WINDOW_EDGE_1 = 3'd2;  // Reading: flux detected, wait half window
    localparam SW_WINDOW_LOAD   = 3'd3;  // Writing: load shift register
    localparam SW_WINDOW_MIDDLE = 3'd4;  // Writing: check MSB
    localparam SW_WINDOW_END    = 3'd5;  // Writing: end window
    localparam SW_UNDERRUN      = 3'd6;  // Writing: underrun error

    reg [2:0]  rw_state;
    reg [5:0]  window_counter; // Countdown for window timing

    //=========================================================================
    // Window Timing (from MAME iwm.cpp half_window_size/window_size)
    //=========================================================================
    // Window timing depends on drive type:
    //
    // IMPORTANT: Window timing runs at 14M for precision!
    // MAME uses cycle counts at 7MHz, but processes flux at exact arrival times.
    // vsim samples at discrete clock edges, so we run at 14M to minimize
    // quantization error. Without 14M precision, flux arrival time is rounded
    // to 7M edges, causing 0-1 cycle error per bit that accumulates and
    // causes byte boundary drift.
    //
    // Window timing in 14M cycles (doubled from MAME's 7MHz values):
    // MAME mode 0x00 (slow): half=14@7M, window=28@7M -> half=28@14M, window=56@14M (4µs)
    // MAME mode 0x08 (fast): half=7@7M, window=14@7M -> half=14@14M, window=28@14M (2µs)
    // Note: 3.5" drives use 2µs bit cells but ROM often doesn't set fast mode bit!

    wire        fast_mode = SW_MODE[3];
    // Window timing: MAME uses 7MHz clock, we run at 14MHz.
    // For 3.5" drives: 2µs bit cells, window = 28 @ 14MHz (matches MAME mode 0x08 fast)
    // For 5.25" drives: 4µs bit cells (slow) or 2µs (fast)
    // Note: ROM typically sets mode=0x0F for 3.5" drives (fast mode + async).
    wire [5:0]  full_window = IS_35_INCH ? 6'd28 : (fast_mode ? 6'd28 : 6'd56);
    wire [5:0]  half_window = IS_35_INCH ? 6'd14 : (fast_mode ? 6'd14 : 6'd28);

    //=========================================================================
    // Flux Edge Detection
    //=========================================================================

    reg        prev_flux;
    reg        prev_sm_active;  // For debug: track state machine activation
    reg        flux_pending;    // Latched when flux arrives during EDGE_1
    reg        flux_seen;       // Latched at 14M when flux edge detected, cleared at 7M
    wire       flux_edge = FLUX_TRANSITION && !prev_flux;

`ifdef SIMULATION
    reg [31:0] debug_cycle;
    reg [31:0] byte_counter;  // Sequential byte counter for comparison with MAME
    reg [31:0] bytes_read_counter;  // How many bytes CPU has read (valid reads with bit7=1)
    reg [31:0] bytes_lost_counter;  // How many bytes were cleared by async_update before CPU read
`endif

    //=========================================================================
    // State Machine and Data Register Logic
    //=========================================================================

    always @(posedge CLK_14M or posedge RESET) begin
        if (RESET) begin
            rw_state       <= S_IDLE;
            m_rsh          <= 8'h00;
            m_data         <= 8'h00;
            m_whd          <= 8'hBF;  // MAME: initialized to 0xBF
            async_update   <= 4'd0;
            bit7_acknowledged <= 1'b0;
            m_data_read    <= 1'b1;   // Start as "read" so first byte triggers ready
            m_rw_mode      <= 1'b0;   // Start in read mode
            m_motor_was_on <= 1'b0;
            window_counter <= 6'd0;
            prev_flux      <= 1'b0;
            prev_sm_active <= 1'b0;
            flux_pending   <= 1'b0;
            flux_seen      <= 1'b0;
            rd_latched     <= 1'b0;
`ifdef SIMULATION
            debug_cycle    <= 32'd0;
            byte_counter   <= 32'd0;
            bytes_read_counter <= 32'd0;
            bytes_lost_counter <= 32'd0;
`endif
        end else begin
`ifdef SIMULATION
            debug_cycle <= debug_cycle + 1;
`endif
            // MAME behavior: Clear m_data when entering read mode
            // Only reset if motor was truly stopped (not spinning), not just command toggling
            if (MOTOR_ACTIVE && !m_motor_was_on && !SW_Q7 && !MOTOR_SPINNING) begin
                m_data <= 8'h00;
                m_rw_mode <= 1'b0;
                rw_state <= S_IDLE;
`ifdef SIMULATION
                $display("IWM_FLUX: Entering READ mode, m_data <= 0x00");
`endif
            end else if (MOTOR_ACTIVE && m_motor_was_on && m_rw_mode && !SW_Q7) begin
                // Switching from write mode to read mode - always reset
                m_data <= 8'h00;
                m_rw_mode <= 1'b0;
                rw_state <= S_IDLE;
`ifdef SIMULATION
                $display("IWM_FLUX: Switching to READ mode, m_data <= 0x00");
`endif
            end else if (MOTOR_ACTIVE && SW_Q7 && !m_rw_mode) begin
                m_rw_mode <= 1'b1;
                m_whd <= m_whd | 8'h40;
            end else if (!MOTOR_ACTIVE && m_motor_was_on) begin
                // Motor command off - but only reset state if motor actually stopped
                m_whd <= m_whd & 8'hBF;
                m_rw_mode <= 1'b0;
                // Don't reset state if motor is still spinning - bytes may still be decoding
                if (!MOTOR_SPINNING) begin
                    rw_state <= S_IDLE;
                end
`ifdef SIMULATION
                $display("IWM_FLUX: Motor off, m_whd <= %02h (cleared bit 6) spin=%0d", m_whd & 8'hBF, MOTOR_SPINNING);
`endif
            end
            m_motor_was_on <= MOTOR_ACTIVE;

            // MAME async_update logic - NOTE: Countdown runs at 7MHz (see CLK_7M_EN block below)
            // In async mode, m_data is cleared 14 cycles (at 7MHz, ~2µs) after a valid byte was read.
            // This happens BEFORE the next read is processed, so the read sees 0x00.

            // Always track flux edges at 14M (so we don't miss any)
            prev_flux <= FLUX_TRANSITION;

            // Latch flux edge at 14M for processing at 7M
            if (flux_edge) begin
                flux_seen <= 1'b1;
            end

            // MAME async_update countdown at 7MHz (matches iwm.cpp update_phases logic)
            // After CPU reads valid byte, m_data is cleared after 14 7M-cycles (~2µs)
            if (CLK_7M_EN) begin
                if (async_update != 0) begin
                    if (async_update == 1) begin
                        // Counter about to hit 0 - clear m_data NOW (unless byte completing)
                        if (is_async && !byte_completing) begin
`ifdef SIMULATION
                            // CRITICAL: If m_data_read is still 0, CPU never read this byte!
                            if (!m_data_read && m_data[7]) begin
                                bytes_lost_counter <= bytes_lost_counter + 1;
                                $display("IWM_FLUX: *** BYTE LOST #%0d *** ASYNC_UPDATE_EXPIRED clearing UNREAD m_data=%02h (completed=%0d read=%0d) @cycle=%0d",
                                         bytes_lost_counter + 1, m_data, byte_counter, bytes_read_counter, debug_cycle);
                            end else begin
                                $display("IWM_FLUX: ASYNC_UPDATE_EXPIRED clearing m_data (was %02h, was_read=%0d) @cycle=%0d",
                                         m_data, m_data_read, debug_cycle);
                            end
`endif
                            m_data <= 8'h00;
                            bit7_acknowledged <= 1'b0;
                        end
                    end
                    async_update <= async_update - 1'b1;
                end
            end

            // State machine runs at 14M for precise flux timing!
            // MAME's IWM clocks at 7M but processes flux at exact arrival times.
            // vsim must run at 14M to avoid timing quantization that causes
            // byte boundary drift. Window values are doubled to compensate.
`ifdef SIMULATION
            if ((MOTOR_SPINNING && DISK_READY) != prev_sm_active) begin
                $display("IWM_FLUX: State machine %s (MOTOR_SPINNING=%0d DISK_READY=%0d)",
                         (MOTOR_SPINNING && DISK_READY) ? "ACTIVE" : "IDLE",
                         MOTOR_SPINNING, DISK_READY);
            end
`endif
            if (MOTOR_SPINNING && DISK_READY) begin
                case (rw_state)
                    S_IDLE: begin
                        rw_state <= SR_WINDOW_EDGE_0;
                        window_counter <= full_window;
                        m_rsh <= 8'h00;
                        flux_seen <= 1'b0;  // Clear on state machine start
`ifdef BYTE_FRAME_DEBUG
                        $display("BYTE_START: pos=%0d window=%0d half=%0d mode=%02h",
                                 DISK_BIT_POSITION, full_window, half_window, SW_MODE);
`else
`ifdef SIMULATION
                        $display("IWM_FLUX: START_READ cycle=%0d win=%0d mode=%02h",
                                 debug_cycle, full_window, SW_MODE);
`endif
`endif
                    end

                    SR_WINDOW_EDGE_0: begin
                        // Check for flux edge (latched at 14M) OR pending flux from EDGE_1
                        if (flux_seen || flux_pending) begin
                            rw_state <= SR_WINDOW_EDGE_1;
                            // CRITICAL FIX: Anchor half-window to flux arrival, like MAME
                            // MAME sets m_next_state_change = flux_time + half_window
                            // When flux arrives early in window, we need to wait longer
                            // When flux arrives late, we wait shorter (but at least 1 cycle)
                            // The flux arrived at the current cycle, so half_window from now
                            // is correct. But we also need to account for where we were
                            // in the window when flux arrived.
                            //
                            // For a 28-cycle window with half=14:
                            // - If flux arrives when window_counter=20, we're 8 cycles into window
                            // - Expected flux at cycle 14 (middle), actual at cycle 8
                            // - Wait half_window (14) to reach cycle 22, bit boundary at 28
                            //
                            // Actually, the MAME behavior is simpler: just wait half_window
                            // from flux arrival. The next window then starts fresh.
                            // The key is that consecutive 1-bits work because flux_pending
                            // captures early flux during EDGE_1.
                            window_counter <= half_window;
                            flux_pending <= 1'b0;  // Clear pending flag
                            flux_seen <= 1'b0;     // Clear seen flag after processing
`ifdef BYTE_FRAME_DEBUG
                            $display("BYTE_FLUX: pos=%0d flux_detected win_remain=%0d->half=%0d pending=%0d sr=%02h",
                                     DISK_BIT_POSITION, window_counter, half_window, flux_pending, m_rsh);
`endif
                        end else if (window_counter == 6'd1) begin
`ifdef BYTE_FRAME_DEBUG
                            $display("BYTE_SHIFT: pos=%0d bit=0 sr=%02h->%02h bitnum=%0d",
                                     DISK_BIT_POSITION, m_rsh, {m_rsh[6:0], 1'b0},
                                     (m_rsh[6] ? 1 : (m_rsh[5] ? 2 : (m_rsh[4] ? 3 : (m_rsh[3] ? 4 : (m_rsh[2] ? 5 : (m_rsh[1] ? 6 : (m_rsh[0] ? 7 : 8))))))));
`endif
                            m_rsh <= {m_rsh[6:0], 1'b0};
                            window_counter <= full_window;
                        end else begin
                            window_counter <= window_counter - 1'd1;
                        end
                    end

                    SR_WINDOW_EDGE_1: begin
                        // MAME behavior: In EDGE_1, don't immediately act on flux - but
                        // latch it so we detect it immediately when we go to EDGE_0.
                        // This handles consecutive 1-bits where flux arrives before
                        // the half-window completes.
                        if (flux_seen) begin
                            flux_pending <= 1'b1;  // Latch for use in EDGE_0
                            flux_seen <= 1'b0;     // Clear seen flag
                        end

                        if (window_counter == 6'd1) begin
`ifdef BYTE_FRAME_DEBUG
                            $display("BYTE_SHIFT: pos=%0d bit=1 sr=%02h->%02h bitnum=%0d",
                                     DISK_BIT_POSITION, m_rsh, {m_rsh[6:0], 1'b1},
                                     (m_rsh[6] ? 1 : (m_rsh[5] ? 2 : (m_rsh[4] ? 3 : (m_rsh[3] ? 4 : (m_rsh[2] ? 5 : (m_rsh[1] ? 6 : (m_rsh[0] ? 7 : 8))))))));
`endif
                            m_rsh <= {m_rsh[6:0], 1'b1};
                            rw_state <= SR_WINDOW_EDGE_0;
                            window_counter <= full_window;
                        end else begin
                            window_counter <= window_counter - 1'd1;
                        end
                    end

                    default: begin
                        rw_state <= S_IDLE;
                    end
                endcase

                // Byte complete when MSB is set
                if (m_rsh >= 8'h80) begin
`ifdef SIMULATION
                    byte_counter <= byte_counter + 1;
`endif
`ifdef BYTE_FRAME_DEBUG
                    $display("BYTE_FORMED: pos=%0d byte#=%0d data=%02h",
                             DISK_BIT_POSITION, byte_counter + 1, m_rsh);
`else
`ifdef SIMULATION
                    $display("IWM_FLUX: BYTE_COMPLETE_ASYNC data=%02h pos=%0d byte#=%0d @cycle=%0d",
                             m_rsh, DISK_BIT_POSITION, byte_counter + 1, debug_cycle);
`endif
`endif
                    m_data <= m_rsh;
                    m_rsh <= 8'h00;
                    m_data_read <= 1'b0;
                    // MAME behavior: Reset async_update when new byte completes.
                    // Also clear bit7_acknowledged so the new byte's bit 7 is visible.
                    bit7_acknowledged <= 1'b0;
                    async_update <= 6'd0;
                end
            end

            // Reset state when motor stops or disk removed
            if (!MOTOR_SPINNING || !DISK_READY) begin
                rw_state <= S_IDLE;
                window_counter <= 6'd0;
                flux_pending <= 1'b0;
                flux_seen <= 1'b0;
                bit7_acknowledged <= 1'b0;
                async_update <= 4'd0;
            end

            prev_sm_active <= MOTOR_SPINNING && DISK_READY;

            // CPU read edge detection: clear latch when RD goes low
            if (!RD || !CEN) begin
                if (rd_latched) begin
                    // CPU read just finished - NOW acknowledge bit 7
                    // This ensures the FIRST read sees bit 7=1, but subsequent ones see 0
                    // CRITICAL: Only set if this was a DATA register read (m_data_read was set)
                    // AND a new byte is NOT currently completing!
                    if (MOTOR_ACTIVE && is_async && effective_data_raw[7] && m_data_read && !byte_completing) begin
                        bit7_acknowledged <= 1'b1;
`ifdef SIMULATION
                        $display("IWM_FLUX: BIT7_ACKNOWLEDGED set (data=%02h) @cycle=%0d", effective_data_raw, debug_cycle);
`endif

                        // MAME async mode behavior:
                        // Start countdown to clear the entire byte after 14 cycles (2us).
                        // By starting it here (at the end of the read), we ensure the
                        // data remains valid for the full duration of the CPU access.
                        if (async_update == 0) begin
                            async_update <= 6'd14; // 14 cycles at 7MHz = 2µs (matches MAME)
`ifdef SIMULATION
                            $display("IWM_FLUX: async_update started (14 7M-cycles) @cycle=%0d", debug_cycle);
`endif
                        end
                    end
                end
                rd_latched <= 1'b0;
            end

            // Set data_read flag when CPU reads data register (Q7=0, Q6=0)
            // Use immediate Q6/Q7 values from current address
            // IMPORTANT: Only process ONCE per CPU read cycle using edge detection
            // CEN (phi2) ensures we're in the valid part of the bus cycle
            if (RD && CEN && !rd_latched) begin
                rd_latched <= 1'b1;  // Mark this read as processed
                // Calculate immediate Q6/Q7 inline
                if ((((ADDR[3:1] == 3'b111) ? ADDR[0] : SW_Q7) == 1'b0) &&
                    (((ADDR[3:1] == 3'b110) ? ADDR[0] : SW_Q6) == 1'b0)) begin
                    m_data_read <= 1'b1;
`ifdef SIMULATION
                    // Count valid data reads (bit7=1) for statistics
                    if (MOTOR_ACTIVE && effective_data_raw[7]) begin
                        bytes_read_counter <= bytes_read_counter + 1;
                    end
`endif
                    // Note: async_update now started at END of read (see above)
                end
            end
        end
    end

    //=========================================================================
    // Register Read Logic (Q6/Q7 select)
    //=========================================================================
    // Q7 Q6 | Read Returns
    // ------+-------------
    //  0  0 | Data register (disk byte)
    //  0  1 | Status register
    //  1  0 | Write handshake register
    //  1  1 | 0xFF (or mode bits)

    // Status register (MAME reference: iwm.cpp status_r() line 303)
    // Bit 7: SENSE_BIT - drive status sense line (write-protect, disk present, etc.)
    //        Selected by phase lines, comes from drive via SENSE_BIT input
    // Bit 6: 0 (reserved)
    // Bit 5: motor_active && disk_installed
    // Bits 4-0: mode register
    // Note: data_ready is NOT in the status register - it's only relevant for
    //       determining when to read the DATA register (Q6=0, Q7=0)
    wire motor_status_bit = MOTOR_ACTIVE && DISK_MOUNTED;
    wire [7:0] status_reg = {SENSE_BIT, 1'b0, motor_status_bit, SW_MODE[4:0]};

    // Write handshake register
    wire [7:0] handshake_reg = 8'h80;

    // Immediate Q6/Q7 values for current access
    // If current access is to Q6/Q7 switch, use ADDR[0] for that bit
    // Otherwise use the latched value from SW_Q6/SW_Q7
    wire access_q6 = (ADDR[3:1] == 3'b110);
    wire access_q7 = (ADDR[3:1] == 3'b111);
    wire immediate_q6 = access_q6 ? ADDR[0] : SW_Q6;
    wire immediate_q7 = access_q7 ? ADDR[0] : SW_Q7;

    // Combinatorial bypass for same-cycle read
    // MAME behavior: always return m_data (the completed byte), which holds its value
    // until the next byte completes. The byte_completing bypass handles the case where
    // the CPU reads in the same cycle that m_rsh reaches 0x80+.
    wire byte_completing = (m_rsh >= 8'h80) && MOTOR_SPINNING && DISK_READY;
    wire [7:0] effective_data_raw = byte_completing ? m_rsh : m_data;

    // MAME behavior: mask bit 7 after it has been acknowledged by a CPU read.
    // The bit 7 remains 0 until the next byte completes (clearing bit7_acknowledged).
    // In async mode, the entire byte eventually clears after 14 cycles (2us).
    // CRITICAL: Never mask if a new byte is just completing!
    wire [7:0] effective_data = (MOTOR_ACTIVE && is_async && bit7_acknowledged && !byte_completing) ? 
                                 (effective_data_raw & 8'h7F) : effective_data_raw;

    // Helper wires for byte completion logic to avoid race conditions
    wire cpu_reading_data = RD && !immediate_q7 && !immediate_q6;
    wire cpu_reading_valid_data = cpu_reading_data && MOTOR_ACTIVE && is_async && effective_data_raw[7];

    reg [7:0] data_out_mux;
    always @(*) begin
        case ({immediate_q7, immediate_q6})
            2'b00: data_out_mux = MOTOR_ACTIVE ? effective_data : 8'hFF;
            2'b01: data_out_mux = status_reg;
            2'b10: data_out_mux = handshake_reg;
            2'b11: data_out_mux = 8'hFF;
        endcase
    end

    //=========================================================================
    // Output Assignments
    //=========================================================================

    assign DATA_OUT     = data_out_mux;
    assign FLUX_WRITE   = 1'b0;  // TODO: implement write support
    assign DEBUG_RSH    = m_rsh;
    assign DEBUG_STATE  = rw_state;

`ifdef SIMULATION
    // Debug: log register reads (only on CEN/PH2 to log once per CPU access)
    always @(posedge CLK_14M) begin
        if (RD && CEN) begin
            case ({immediate_q7, immediate_q6})
                2'b00: $display("IWM_FLUX: READ DATA @%01h -> %02h pos=%0d (motor=%0d rsh=%02h data=%02h bc=%0d dr=%0d q6=%0d q7=%0d)",
                               ADDR, data_out_mux, DISK_BIT_POSITION, MOTOR_ACTIVE, m_rsh, m_data, byte_completing, DISK_READY, SW_Q6, SW_Q7);
                2'b01: $display("IWM_FLUX: READ STATUS @%01h -> %02h (sense=%0d m_reg=%01h latched=%01h sel=%0d phases=%04b is_35=%0d motor_active=%0d mounted=%0d)",
                               ADDR, data_out_mux, SENSE_BIT, {DISKREG_SEL, LATCHED_SENSE_REG}, LATCHED_SENSE_REG, DISKREG_SEL, SW_PHASES, IS_35_INCH, MOTOR_ACTIVE, DISK_MOUNTED);
                2'b10: $display("IWM_FLUX: READ HANDSHAKE @%01h -> %02h", ADDR, data_out_mux);
                2'b11: $display("IWM_FLUX: READ @%01h -> %02h (q7=q6=1)", ADDR, data_out_mux);
            endcase
        end

        // Periodic statistics - every 10M cycles (~0.7 seconds)
        if (debug_cycle[23:0] == 24'h0 && debug_cycle > 0 && MOTOR_ACTIVE) begin
            $display("IWM_FLUX: *** STATS @cycle=%0d *** bytes_completed=%0d bytes_read=%0d bytes_lost=%0d loss_rate=%0d%%",
                     debug_cycle, byte_counter, bytes_read_counter, bytes_lost_counter,
                     (byte_counter > 0) ? (bytes_lost_counter * 100 / byte_counter) : 0);
        end
    end
`endif

    //=========================================================================
    // Sector Read Tracking (for debug - tracks byte stream, not CPU reads)
    //=========================================================================
    // This state machine watches the byte stream (m_data) and tracks sector reads.
    // 3.5" GCR format:
    //   Address field: D5 AA 96 <track> <sector> <side> <format> <checksum> DE AA
    //   Data field:    D5 AA AD <12 tag> <512 data> <4 checksum> DE AA
    // Note: This tracks raw bytes from the disk, independent of CPU read timing.

`ifdef SECTOR_DEBUG
    // GCR 6-2 decode function for 3.5" disk address fields
    // Input: raw GCR byte (0x80-0xFF), Output: decoded 6-bit value (0x00-0x3F, or 0x80 for invalid)
    // Table from Clemens emulator (clem_disk.c)
    function [7:0] gcr_6_2_decode;
        input [7:0] gcr_byte;
        begin
            case (gcr_byte)
                // 0x90-0x97
                8'h96: gcr_6_2_decode = 8'h00;
                8'h97: gcr_6_2_decode = 8'h01;
                // 0x98-0x9F
                8'h9A: gcr_6_2_decode = 8'h02;
                8'h9B: gcr_6_2_decode = 8'h03;
                8'h9D: gcr_6_2_decode = 8'h04;
                8'h9E: gcr_6_2_decode = 8'h05;
                8'h9F: gcr_6_2_decode = 8'h06;
                // 0xA0-0xA7
                8'hA6: gcr_6_2_decode = 8'h07;
                8'hA7: gcr_6_2_decode = 8'h08;
                // 0xA8-0xAF
                8'hAB: gcr_6_2_decode = 8'h09;
                8'hAC: gcr_6_2_decode = 8'h0A;
                8'hAD: gcr_6_2_decode = 8'h0B;
                8'hAE: gcr_6_2_decode = 8'h0C;
                8'hAF: gcr_6_2_decode = 8'h0D;
                // 0xB0-0xB7
                8'hB2: gcr_6_2_decode = 8'h0E;
                8'hB3: gcr_6_2_decode = 8'h0F;
                8'hB4: gcr_6_2_decode = 8'h10;
                8'hB5: gcr_6_2_decode = 8'h11;
                8'hB6: gcr_6_2_decode = 8'h12;
                8'hB7: gcr_6_2_decode = 8'h13;
                // 0xB8-0xBF
                8'hB9: gcr_6_2_decode = 8'h14;
                8'hBA: gcr_6_2_decode = 8'h15;
                8'hBB: gcr_6_2_decode = 8'h16;
                8'hBC: gcr_6_2_decode = 8'h17;
                8'hBD: gcr_6_2_decode = 8'h18;
                8'hBE: gcr_6_2_decode = 8'h19;
                8'hBF: gcr_6_2_decode = 8'h1A;
                // 0xC8-0xCF
                8'hCB: gcr_6_2_decode = 8'h1B;
                8'hCD: gcr_6_2_decode = 8'h1C;
                8'hCE: gcr_6_2_decode = 8'h1D;
                8'hCF: gcr_6_2_decode = 8'h1E;
                // 0xD0-0xD7
                8'hD3: gcr_6_2_decode = 8'h1F;
                8'hD6: gcr_6_2_decode = 8'h20;
                8'hD7: gcr_6_2_decode = 8'h21;
                // 0xD8-0xDF
                8'hD9: gcr_6_2_decode = 8'h22;
                8'hDA: gcr_6_2_decode = 8'h23;
                8'hDB: gcr_6_2_decode = 8'h24;
                8'hDC: gcr_6_2_decode = 8'h25;
                8'hDD: gcr_6_2_decode = 8'h26;
                8'hDE: gcr_6_2_decode = 8'h27;
                8'hDF: gcr_6_2_decode = 8'h28;
                // 0xE0-0xE7
                8'hE5: gcr_6_2_decode = 8'h29;
                8'hE6: gcr_6_2_decode = 8'h2A;
                8'hE7: gcr_6_2_decode = 8'h2B;
                // 0xE8-0xEF
                8'hE9: gcr_6_2_decode = 8'h2C;
                8'hEA: gcr_6_2_decode = 8'h2D;
                8'hEB: gcr_6_2_decode = 8'h2E;
                8'hEC: gcr_6_2_decode = 8'h2F;
                8'hED: gcr_6_2_decode = 8'h30;
                8'hEE: gcr_6_2_decode = 8'h31;
                8'hEF: gcr_6_2_decode = 8'h32;
                // 0xF0-0xF7
                8'hF2: gcr_6_2_decode = 8'h33;
                8'hF3: gcr_6_2_decode = 8'h34;
                8'hF4: gcr_6_2_decode = 8'h35;
                8'hF5: gcr_6_2_decode = 8'h36;
                8'hF6: gcr_6_2_decode = 8'h37;
                8'hF7: gcr_6_2_decode = 8'h38;
                // 0xF8-0xFF
                8'hF9: gcr_6_2_decode = 8'h39;
                8'hFA: gcr_6_2_decode = 8'h3A;
                8'hFB: gcr_6_2_decode = 8'h3B;
                8'hFC: gcr_6_2_decode = 8'h3C;
                8'hFD: gcr_6_2_decode = 8'h3D;
                8'hFE: gcr_6_2_decode = 8'h3E;
                8'hFF: gcr_6_2_decode = 8'h3F;
                default: gcr_6_2_decode = 8'h80;  // Invalid GCR byte
            endcase
        end
    endfunction

    // Sector tracking state machine
    localparam SEC_IDLE       = 4'd0;
    localparam SEC_WAIT_AA1   = 4'd1;  // Saw D5, waiting for first AA
    localparam SEC_WAIT_96    = 4'd2;  // Saw D5 AA, waiting for 96 (addr) or AD (data)
    localparam SEC_ADDR_TRACK = 4'd3;  // Reading address field: track byte
    localparam SEC_ADDR_SEC   = 4'd4;  // Reading address field: sector byte
    localparam SEC_ADDR_SIDE  = 4'd5;  // Reading address field: side byte
    localparam SEC_ADDR_FMT   = 4'd6;  // Reading address field: format byte
    localparam SEC_ADDR_CSUM  = 4'd7;  // Reading address field: checksum byte
    localparam SEC_DATA_TAG   = 4'd8;  // Reading data field: 12 tag bytes
    localparam SEC_DATA_READ  = 4'd9;  // Reading data field: 512 data bytes
    localparam SEC_DATA_CSUM  = 4'd10; // Reading data field: 4 checksum bytes

    reg [3:0]  sec_state;
    reg [7:0]  sec_track;         // Raw GCR byte
    reg [7:0]  sec_sector;        // Raw GCR byte
    reg [7:0]  sec_side;          // Raw GCR byte
    reg [7:0]  sec_format;        // Raw GCR byte
    reg [7:0]  sec_addr_csum;     // Raw checksum byte from address field
    reg [5:0]  sec_decoded_track; // Decoded 6-bit track value
    reg [5:0]  sec_decoded_sector;// Decoded 6-bit sector value
    reg [5:0]  sec_decoded_side;  // Decoded 6-bit side value
    reg [5:0]  sec_decoded_format;// Decoded 6-bit format value
    reg [5:0]  sec_running_xor;   // Running XOR of decoded values (should be 0 after all 5 bytes)
    reg [9:0]  sec_data_count;    // Counter for data bytes (0-511)
    reg [3:0]  sec_tag_count;     // Counter for tag bytes (0-11)
    reg [1:0]  sec_csum_count;    // Counter for checksum bytes (0-3)
    reg [31:0] sec_data_csum;     // Running checksum for data field (3 bytes used)
    reg [16:0] sec_start_pos;     // Position where sector started (for logging)

    // Statistics
    reg [15:0] sec_addr_ok_count;
    reg [15:0] sec_addr_fail_count;
    reg [15:0] sec_data_count_total;

    // Detect byte completion using m_rsh >= 0x80 signal (byte_completing is defined earlier)
    // Use edge detection since byte_completing is a level signal during the completion cycle.
    reg        prev_byte_completing;
    wire       new_byte = byte_completing && !prev_byte_completing;

    always @(posedge CLK_14M or posedge RESET) begin
        if (RESET) begin
            sec_state <= SEC_IDLE;
            sec_track <= 8'd0;
            sec_sector <= 8'd0;
            sec_side <= 8'd0;
            sec_format <= 8'd0;
            sec_addr_csum <= 8'd0;
            sec_decoded_track <= 6'd0;
            sec_decoded_sector <= 6'd0;
            sec_decoded_side <= 6'd0;
            sec_decoded_format <= 6'd0;
            sec_running_xor <= 6'd0;
            sec_data_count <= 10'd0;
            sec_tag_count <= 4'd0;
            sec_csum_count <= 2'd0;
            sec_data_csum <= 32'd0;
            sec_start_pos <= 17'd0;
            sec_addr_ok_count <= 16'd0;
            sec_addr_fail_count <= 16'd0;
            sec_data_count_total <= 16'd0;
            prev_byte_completing <= 1'b0;
        end else if (MOTOR_SPINNING && DISK_READY) begin
            prev_byte_completing <= byte_completing;

            // State machine triggered by new bytes
            // NOTE: When new_byte fires (byte_completing edge), the completed byte is in m_rsh
            if (new_byte) begin
                case (sec_state)
                    SEC_IDLE: begin
                        if (m_rsh == 8'hD5) begin
                            sec_state <= SEC_WAIT_AA1;
                            sec_start_pos <= DISK_BIT_POSITION;
                        end
                    end

                    SEC_WAIT_AA1: begin
                        if (m_rsh == 8'hAA)
                            sec_state <= SEC_WAIT_96;
                        else if (m_rsh == 8'hD5)
                            sec_state <= SEC_WAIT_AA1;  // Stay, could be new marker
                        else
                            sec_state <= SEC_IDLE;
                    end

                    SEC_WAIT_96: begin
                        if (m_rsh == 8'h96) begin
                            // Address field prologue complete
                            sec_state <= SEC_ADDR_TRACK;
                            $display("SECTOR: D5 AA 96 at pos=%0d (address prologue)", sec_start_pos);
                        end else if (m_rsh == 8'hAD) begin
                            // Data field prologue
                            sec_state <= SEC_DATA_TAG;
                            sec_tag_count <= 4'd0;
                            $display("SECTOR: D5 AA AD at pos=%0d (data prologue) for T%0d S%0d",
                                     sec_start_pos, sec_track, sec_sector);
                        end else if (m_rsh == 8'hD5) begin
                            sec_state <= SEC_WAIT_AA1;
                            sec_start_pos <= DISK_BIT_POSITION;
                        end else begin
                            sec_state <= SEC_IDLE;
                        end
                    end

                    SEC_ADDR_TRACK: begin
                        sec_track <= m_rsh;
                        sec_decoded_track <= gcr_6_2_decode(m_rsh)[5:0];
                        sec_running_xor <= gcr_6_2_decode(m_rsh)[5:0];  // Start running XOR
                        sec_state <= SEC_ADDR_SEC;
                    end

                    SEC_ADDR_SEC: begin
                        sec_sector <= m_rsh;
                        sec_decoded_sector <= gcr_6_2_decode(m_rsh)[5:0];
                        sec_running_xor <= sec_running_xor ^ gcr_6_2_decode(m_rsh)[5:0];
                        sec_state <= SEC_ADDR_SIDE;
                    end

                    SEC_ADDR_SIDE: begin
                        sec_side <= m_rsh;
                        sec_decoded_side <= gcr_6_2_decode(m_rsh)[5:0];
                        sec_running_xor <= sec_running_xor ^ gcr_6_2_decode(m_rsh)[5:0];
                        sec_state <= SEC_ADDR_FMT;
                    end

                    SEC_ADDR_FMT: begin
                        sec_format <= m_rsh;
                        sec_decoded_format <= gcr_6_2_decode(m_rsh)[5:0];
                        sec_running_xor <= sec_running_xor ^ gcr_6_2_decode(m_rsh)[5:0];
                        sec_state <= SEC_ADDR_CSUM;
                    end

                    SEC_ADDR_CSUM: begin
                        sec_addr_csum <= m_rsh;
                        // ROM-style validation: XOR of all 5 decoded bytes must equal 0
                        // The checksum byte is chosen so that track^sector^side^format^checksum = 0
                        if ((sec_running_xor ^ gcr_6_2_decode(m_rsh)[5:0]) == 6'd0) begin
                            sec_addr_ok_count <= sec_addr_ok_count + 1;
                            $display("SECTOR: ADDR OK T=%0d S=%0d side=%02h fmt=%02h (raw: %02h %02h %02h %02h %02h) pos=%0d",
                                     sec_decoded_track, sec_decoded_sector, sec_decoded_side, sec_decoded_format,
                                     sec_track, sec_sector, sec_side, sec_format, m_rsh, DISK_BIT_POSITION);
                        end else begin
                            sec_addr_fail_count <= sec_addr_fail_count + 1;
                            $display("SECTOR: ADDR FAIL T=%0d S=%0d side=%02h fmt=%02h xor=%02h (raw: %02h %02h %02h %02h %02h) pos=%0d",
                                     sec_decoded_track, sec_decoded_sector, sec_decoded_side, sec_decoded_format,
                                     sec_running_xor ^ gcr_6_2_decode(m_rsh)[5:0],
                                     sec_track, sec_sector, sec_side, sec_format, m_rsh, DISK_BIT_POSITION);
                        end
                        sec_state <= SEC_IDLE;  // Wait for data field
                    end

                    SEC_DATA_TAG: begin
                        sec_tag_count <= sec_tag_count + 1;
                        if (sec_tag_count == 4'd11) begin
                            sec_state <= SEC_DATA_READ;
                            sec_data_count <= 10'd0;
                            sec_data_csum <= 32'd0;
                        end
                    end

                    SEC_DATA_READ: begin
                        // Track data bytes (simplified - not computing full checksum)
                        sec_data_count <= sec_data_count + 1;
                        if (sec_data_count == 10'd511) begin
                            sec_state <= SEC_DATA_CSUM;
                            sec_csum_count <= 2'd0;
                            sec_data_count_total <= sec_data_count_total + 1;
                        end
                    end

                    SEC_DATA_CSUM: begin
                        sec_csum_count <= sec_csum_count + 1;
                        if (sec_csum_count == 2'd3) begin
                            $display("SECTOR: DATA COMPLETE T=%02h S=%02h (512 bytes read) pos=%0d",
                                     sec_track, sec_sector, DISK_BIT_POSITION);
                            sec_state <= SEC_IDLE;
                        end
                    end

                    default: sec_state <= SEC_IDLE;
                endcase
            end

            // Reset if marker sequence broken
            if (!MOTOR_SPINNING || !DISK_READY) begin
                sec_state <= SEC_IDLE;
            end
        end
    end

    // Periodic statistics for sector tracking
    always @(posedge CLK_14M) begin
        if (debug_cycle[24:0] == 25'h0 && debug_cycle > 0 && MOTOR_ACTIVE) begin
            $display("SECTOR: *** STATS *** addr_ok=%0d addr_fail=%0d data_complete=%0d",
                     sec_addr_ok_count, sec_addr_fail_count, sec_data_count_total);
        end
    end
`endif

endmodule
