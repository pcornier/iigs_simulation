
module mcode(CLK, RST_N, EN, IR, STATE, M);
   input       CLK;
   input       RST_N;
   input       EN;
   input [7:0] IR;
   input [3:0] STATE;
   output MCode_r   M;

parameter [51:0] M_TAB[0:2047] = '{
{3'b111, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b100, 2'b10},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b010, 2'b10},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b010, 2'b10},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b001, 2'b10},
{3'b000, 3'b100, 2'b00, 3'b010, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b10, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b100, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b010, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b111, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b100, 2'b10},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b010, 2'b10},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b010, 2'b10},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b001, 2'b10},
{3'b000, 3'b100, 2'b00, 3'b010, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b10, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b100, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b010, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 3'b011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01111, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 3'b011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01010, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b10, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b001, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b100, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b01},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b01},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000010, 5'b01010, 2'b11, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b011000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b011000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b110, 3'b001, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b001, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b001, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01111, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b110, 3'b001, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b001, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b001, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01010, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b011, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b100, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b001, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 3'b011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01110, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 3'b011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01010, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b10, 3'b000, 2'b00, 2'b01, 8'b00000101, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b100, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 3'b000, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000010, 5'b00011, 2'b11, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b100, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b110, 3'b001, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b001, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b001, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01110, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 3'b101, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b101, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b101, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01010, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000101, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00100, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00100, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b010, 2'b10},
{3'b010, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b110, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b010, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b100, 2'b10},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b10, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b010, 2'b10},
{3'b010, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b110, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b010, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b01001, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b01001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 3'b011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01100, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b10, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 3'b010, 2'b00, 3'b011, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b100, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b01},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b01},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000010, 5'b01100, 2'b11, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b010, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b01, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b01001, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b01001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b110, 3'b001, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b001, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b001, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01100, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b011, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b100, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b001, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b01001, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b01001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 3'b011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01100, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b10, 3'b000, 2'b00, 2'b01, 8'b00000101, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b100, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 3'b000, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000010, 5'b00010, 2'b11, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b101010, 5'b00001, 2'b11, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b01001, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b01001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 3'b101, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b101, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b101, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01100, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000101, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00101, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00101, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b010, 2'b00, 3'b011, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b111, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b010, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b10, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b11, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b10, 8'b00000001, 3'b001, 3'b000, 3'b110, 2'b00, 6'b001010, 5'b00010, 2'b11, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b11, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b010010, 5'b00010, 2'b11, 3'b000, 2'b10},
{3'b000, 3'b001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b110, 2'b10},
{3'b000, 3'b001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b111, 3'b000, 3'b101, 2'b00, 6'b000101, 5'b10000, 2'b11, 3'b000, 2'b00},
{3'b010, 3'b001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 3'b011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01011, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b10, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b110, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b001, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b001, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b100, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b01},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b01},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000010, 5'b01011, 2'b11, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b110000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b010, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b110, 3'b001, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b001, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b001, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01011, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b011, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b100, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b001, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b11, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b10, 8'b00000001, 3'b001, 3'b000, 3'b110, 2'b00, 6'b001010, 5'b00011, 2'b11, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b11, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b010010, 5'b00011, 2'b11, 3'b000, 2'b10},
{3'b000, 3'b001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b110, 2'b10},
{3'b000, 3'b001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b111, 3'b000, 3'b101, 2'b00, 6'b000101, 5'b10000, 2'b11, 3'b000, 2'b00},
{3'b010, 3'b001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 3'b011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01011, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b10, 3'b000, 2'b00, 2'b01, 8'b00000101, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b100, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 3'b000, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b110, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b011, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b011, 2'b00, 6'b010000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b011, 2'b00, 6'b010000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b01, 6'b000010, 5'b00001, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b110, 3'b000, 3'b000, 2'b10, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 3'b101, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b101, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b101, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01011, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000101, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00110, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00110, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b010, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b010, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01101100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b011, 2'b10},
{3'b010, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b011, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b111, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b111, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 3'b011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01101, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b10, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b010, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b010, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b010, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b100, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b01},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b01},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000010, 5'b01101, 2'b11, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b010, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b010, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b10, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b110, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b010, 3'b110, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b010, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b110, 3'b001, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b001, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b001, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01101, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b011, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b100, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b001, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b111, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b111, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 3'b011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01101, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b10, 3'b000, 2'b00, 2'b01, 8'b00000101, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b100, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 3'b000, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b010, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b010, 3'b111, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b010, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b011010, 5'b00001, 2'b11, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b111, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b010, 3'b111, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b010, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 3'b101, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b101, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b101, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000100, 5'b01101, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000101, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00111, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00111, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b011, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b100, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01101100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b011, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b011, 2'b00, 6'b010010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b011, 2'b00, 6'b010010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b010, 2'b00, 6'b001010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b010, 2'b00, 6'b001010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b10, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b010010, 5'b00010, 2'b11, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b100, 3'b000, 2'b00, 3'b111, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b01001, 2'b01, 3'b000, 2'b01},
{3'b010, 3'b000, 2'b00, 3'b111, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b01001, 2'b10, 3'b000, 2'b01},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b001010, 5'b00000, 2'b11, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b111010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b011, 2'b00, 6'b010010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b011, 2'b00, 6'b010010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b010, 2'b00, 6'b001010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b010, 2'b00, 6'b001010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b011, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b100, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00100, 2'b01, 3'b101, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b011, 2'b00, 6'b010010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b011, 2'b00, 6'b010010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b01, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b010, 2'b00, 6'b001010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b010, 2'b00, 6'b001010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b10, 3'b000, 2'b00, 2'b01, 8'b00000101, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b010010, 5'b00000, 2'b11, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b101, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b001010, 5'b00000, 2'b11, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b111, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b111, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b111, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b111, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000101, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b100, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b111, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b01},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b111, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b01},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b100, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b110, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b01},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b110, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b01},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b10, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b000010, 5'b00000, 2'b11, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b100, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b01},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b01},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b000010, 5'b00000, 2'b11, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 3'b010, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b11, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b011, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b100, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b001, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b01, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b10, 3'b000, 2'b00, 2'b01, 8'b00000101, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b100, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 3'b000, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b101010, 5'b00001, 2'b11, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b010010, 5'b00000, 2'b11, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 3'b000, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000101, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b100, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b011, 2'b00, 6'b010000, 5'b10000, 2'b01, 3'b000, 2'b01},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b011, 2'b00, 6'b010001, 5'b10000, 2'b10, 3'b000, 2'b01},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b010, 3'b000, 2'b00, 3'b110, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b011, 2'b00, 6'b010000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b011, 2'b00, 6'b010001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 3'b011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100010, 5'b00010, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b10, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b111, 2'b00, 6'b010010, 5'b00011, 2'b11, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b100, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b01},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b01},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b001010, 5'b00010, 2'b11, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b011, 2'b00, 6'b010000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b011, 2'b00, 6'b010001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b110, 3'b001, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b001, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b001, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100010, 5'b00010, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b011, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b100, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b001, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b011, 2'b10},
{3'b010, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b011, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 3'b011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100010, 5'b00010, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b10, 3'b000, 2'b00, 2'b01, 8'b00000101, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b100, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 3'b000, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b110, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b010, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b010, 2'b00, 6'b001000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b010, 2'b00, 6'b001000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b110, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b110, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b010, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b010, 3'b110, 2'b10, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b10, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 3'b101, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b101, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b101, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100010, 5'b00010, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000101, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b100, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b010, 2'b00, 6'b001000, 5'b10000, 2'b01, 3'b000, 2'b01},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b010, 2'b00, 6'b001001, 5'b10000, 2'b10, 3'b000, 2'b01},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b010, 3'b000, 2'b00, 3'b110, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b010, 2'b00, 6'b001000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b010, 2'b00, 6'b001001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 3'b011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100010, 5'b00011, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b10, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b001010, 5'b00011, 2'b11, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b100, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b01},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b01},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b00000, 2'b11, 3'b000, 2'b00},
{3'b010, 3'b000, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b001, 2'b00, 6'b000010, 5'b00000, 2'b01, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b010, 2'b00, 6'b001000, 5'b10000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b010, 2'b00, 6'b001001, 5'b10000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b110, 3'b001, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b001, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b001, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100010, 5'b00011, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b001, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b001, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000001, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b011, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b100, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b010, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b001, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b001, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b001, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110111, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00001000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b011, 2'b10},
{3'b010, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b011, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b011, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b011, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10010000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 3'b011, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b011, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100010, 5'b00011, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b101, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b10110100, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00011000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b011, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b01, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b000, 3'b011, 2'b10, 3'b000, 2'b00, 2'b01, 8'b00000101, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b10},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b100, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 3'b000, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b01, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b001, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b010, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b010, 3'b110, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b010, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b110, 2'b00, 6'b000001, 5'b00001, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b010, 3'b000, 2'b00, 3'b101, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b010, 2'b10},
{3'b000, 3'b010, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b011, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b010, 2'b10},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b000, 3'b111, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b010, 3'b111, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b010, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b001, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000011, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000100, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b00},
{3'b110, 3'b101, 2'b00, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b01, 3'b000, 2'b10},
{3'b000, 3'b101, 2'b01, 3'b000, 2'b01, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b10, 3'b000, 2'b10},
{3'b110, 3'b101, 2'b01, 3'b001, 2'b10, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100010, 5'b00011, 2'b11, 3'b000, 2'b00},
{3'b000, 3'b101, 2'b01, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b10, 3'b101, 2'b10},
{3'b010, 3'b101, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b000, 2'b00, 6'b100000, 5'b00000, 2'b01, 3'b101, 2'b10},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b01000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00101000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000101, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b01},
{3'b100, 3'b101, 2'b00, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000000, 5'b01000, 2'b01, 3'b000, 2'b10},
{3'b010, 3'b101, 2'b01, 3'b001, 2'b00, 2'b00, 8'b00000000, 3'b000, 3'b000, 3'b101, 2'b00, 6'b000001, 5'b01000, 2'b10, 3'b000, 2'b10},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX},
{3'bXXX, 3'bXXX, 2'bXX, 3'bXXX, 2'bXX, 2'bXX, 8'bXXXXXXXX, 3'bXXX, 3'bXXX, 3'bXXX, 2'bXX, 6'bXXXXXX, 5'bXXXXX, 2'bXX, 3'bXXX, 2'bXX}};

   parameter [7:0] ALU_TAB[0:16] = '{
      {3'b100, 3'b100, 1'b0, 1'b0},
      {3'b100, 3'b100, 1'b0, 1'b1},
      {3'b110, 3'b100, 1'b0, 1'b0},
      {3'b111, 3'b100, 1'b0, 1'b0},
      {3'b100, 3'b000, 1'b0, 1'b0},
      {3'b100, 3'b001, 1'b0, 1'b0},
      {3'b100, 3'b010, 1'b0, 1'b0},
      {3'b100, 3'b011, 1'b0, 1'b0},
      {3'b100, 3'b111, 1'b1, 1'b0},
      {3'b100, 3'b001, 1'b1, 1'b0},
      {3'b000, 3'b100, 1'b0, 1'b0},
      {3'b010, 3'b100, 1'b0, 1'b0},
      {3'b001, 3'b100, 1'b0, 1'b0},
      {3'b011, 3'b100, 1'b0, 1'b0},
      {3'b100, 3'b101, 1'b0, 1'b0},
      {3'b100, 3'b101, 1'b1, 1'b0},
      {3'b100, 3'b110, 1'b0, 1'b0}
   };

   MicroInst_r         MI;
   ALUCtrl_r        ALUFlags;

   assign ALUFlags = ALU_TAB[MI.ALUCtrl];


   always @(posedge CLK or negedge RST_N)
   begin: xhdl0
      reg [3:0]   STATE2;
      if (RST_N == 1'b0)
         MI <= {3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b11};
      else
      begin
         STATE2 = STATE - 1;
         if (EN == 1'b1)
         begin
            if (STATE == 4'b0000)
               MI <= {3'b000, 3'b000, 2'b00, 3'b000, 2'b00, 2'b00, 8'b00000000, 3'b001, 3'b000, 3'b000, 2'b00, 6'b000000, 5'b00000, 2'b00, 3'b000, 2'b11};
            else
               MI <= M_TAB[({IR, STATE2[2:0]})];
         end
      end
   end

   assign M = {ALUFlags, MI.stateCtrl, MI.addrBus, MI.addrInc, MI.muxCtrl, MI.addrCtrl, MI.loadPC, MI.loadSP, MI.regAXY, MI.loadP, MI.loadT, MI.loadDKB, MI.busCtrl, MI.byteSel, MI.outBus, MI.va};

endmodule
